--
-- This file is automatically generated.  Editing is useless!
--

library ieee;
use ieee.std_logic_1164.all;
use work.fnet_util_pkg.all;

package text_config_data is

  constant text_config_data_size : integer := 2**8;

  type text_config_array_type is array(0 to text_config_data_size-1) of
    std_logic_vector(15 downto 0);

  constant tcfg_index_fixed_ip : integer := 1;
  constant tcfg_index_mac : integer := 2;
  constant tcfg_index_control_ip : integer := 3;
  constant tcfg_index_control_mask : integer := 4;
  constant tcfg_index_int1 : integer := 5;

constant text_config_array : text_config_array_type := (
    i2slv16(16#00c3#), -- [x00] 0x00c3 (x04  3) Branch:  c
    i2slv16(16#0486#), -- [x01] 0x0486 (x13  6) Branch:  f
    i2slv16(16#0689#), -- [x02] 0x0689 (x1b  9) Branch:  i
    i2slv16(16#878d#), -- [x03] 0x878d (x1f 13) Branch:  m
    i2slv16(16#810f#), -- [x04] 0x810f (x05 15) Branch:   o
    i2slv16(16#814e#), -- [x05] 0x814e (x06 14) Branch:    n
    i2slv16(16#8194#), -- [x06] 0x8194 (x07 20) Branch:     t
    i2slv16(16#81d2#), -- [x07] 0x81d2 (x08 18) Branch:      r
    i2slv16(16#820f#), -- [x08] 0x820f (x09 15) Branch:       o
    i2slv16(16#824c#), -- [x09] 0x824c (x0a 12) Branch:        l
    i2slv16(16#829f#), -- [x0a] 0x829f (x0b 31) Branch:         _
    i2slv16(16#0309#), -- [x0b] 0x0309 (x0d  9) Branch:          i
    i2slv16(16#838d#), -- [x0c] 0x838d (x0f 13) Branch:          m
    i2slv16(16#8350#), -- [x0d] 0x8350 (x0e 16) Branch:           p
    i2slv16(16#80f9#), -- [x0e] 0x80f9 (  3  9)  Option:           control_ip
    i2slv16(16#83c1#), -- [x0f] 0x83c1 (x10  1) Branch:           a
    i2slv16(16#8413#), -- [x10] 0x8413 (x11 19) Branch:            s
    i2slv16(16#844b#), -- [x11] 0x844b (x12 11) Branch:            k
    i2slv16(16#8139#), -- [x12] 0x8139 (  4  9)  Option:           control_mask
    i2slv16(16#84c9#), -- [x13] 0x84c9 (x14  9) Branch:   i
    i2slv16(16#8518#), -- [x14] 0x8518 (x15 24) Branch:    x
    i2slv16(16#8545#), -- [x15] 0x8545 (x16  5) Branch:     e
    i2slv16(16#8584#), -- [x16] 0x8584 (x17  4) Branch:      d
    i2slv16(16#85df#), -- [x17] 0x85df (x18 31) Branch:       _
    i2slv16(16#8609#), -- [x18] 0x8609 (x19  9) Branch:        i
    i2slv16(16#8650#), -- [x19] 0x8650 (x1a 16) Branch:         p
    i2slv16(16#8079#), -- [x1a] 0x8079 (  1  9)  Option:         fixed_ip
    i2slv16(16#86ce#), -- [x1b] 0x86ce (x1c 14) Branch:   n
    i2slv16(16#8714#), -- [x1c] 0x8714 (x1d 20) Branch:    t
    i2slv16(16#8761#), -- [x1d] 0x8761 (x1e 33) Branch:     1
    i2slv16(16#8171#), -- [x1e] 0x8171 (  5  1)  Option:     int1
    i2slv16(16#87c1#), -- [x1f] 0x87c1 (x20  1) Branch:   a
    i2slv16(16#8803#), -- [x20] 0x8803 (x21  3) Branch:    c
    i2slv16(16#80b2#), -- [x21] 0x80b2 (  2  2)  Option:    mac
    --
    others => (others => '0')
    );

end text_config_data;
